`timescale 1ns / 1ps
`default_nettype none

module core #(
    parameter int ADDR_WIDTH = 31,
    parameter int DATA_WIDTH = 31
) (
    input i_clk,
    input i_clk_en,
    input i_rst
);

endmodule
