32'd0: o_read_data = 32'd318832704;
32'd4: o_read_data = 32'd4009787396;
32'd8: o_read_data = 32'd1862287369;
32'd12: o_read_data = 32'd326497551;
32'd16: o_read_data = 32'd587243552;
32'd20: o_read_data = 32'd1736441856;
32'd24: o_read_data = 32'd318833151;
32'd28: o_read_data = 32'd589594880;
32'd32: o_read_data = 32'd589697280;
32'd36: o_read_data = 32'd319030528;
32'd40: o_read_data = 32'd54854656;
32'd44: o_read_data = 32'd1662649600;
32'd48: o_read_data = 32'd2199961856;
32'd52: o_read_data = 32'd52723968;
32'd56: o_read_data = 32'd318832897;
32'd60: o_read_data = 32'd1736441856;
32'd64: o_read_data = 32'd319034368;
32'd68: o_read_data = 32'd4025524220;
32'd72: o_read_data = 32'd1878007806;
32'd76: o_read_data = 32'd318833151;
32'd80: o_read_data = 32'd386203648;
32'd84: o_read_data = 32'd319112450;
32'd88: o_read_data = 32'd589697280;
32'd92: o_read_data = 32'd4025540603;
32'd96: o_read_data = 32'd2199961856;
32'd100: o_read_data = 32'd386203648;
32'd104: o_read_data = 32'd319096066;
32'd108: o_read_data = 32'd318832897;
32'd112: o_read_data = 32'd1878040570;
32'd116: o_read_data = 32'd1214606444;
32'd120: o_read_data = 32'd1864397665;
32'd124: o_read_data = 32'd1768714098;
32'd128: o_read_data = 32'd772407296;
32'd132: o_read_data = 32'd1466458484;
32'd136: o_read_data = 32'd661856358;
32'd140: o_read_data = 32'd1869750370;
32'd144: o_read_data = 32'd1919246699;
32'd148: o_read_data = 32'd1717662580;
32'd152: o_read_data = 32'd1057619968;
default: o_read_data = 32'bX; // Default value
