32'd0: o_read_data = 32'd1073742099;
32'd4: o_read_data = 32'd75497711;
32'd8: o_read_data = 32'd155189359;
32'd12: o_read_data = 32'd267744531;
32'd16: o_read_data = 32'd547356707;
32'd20: o_read_data = 32'd32871;
32'd24: o_read_data = 32'd4278255891;
32'd28: o_read_data = 32'd8463395;
32'd32: o_read_data = 32'd1123875;
32'd36: o_read_data = 32'd328723;
32'd40: o_read_data = 32'd279811;
32'd44: o_read_data = 32'd334435;
32'd48: o_read_data = 32'd12656771;
32'd52: o_read_data = 32'd8463363;
32'd56: o_read_data = 32'd16843027;
32'd60: o_read_data = 32'd32871;
32'd64: o_read_data = 32'd1311763;
32'd68: o_read_data = 32'd4238340335;
32'd72: o_read_data = 32'd4263506031;
32'd76: o_read_data = 32'd4278255891;
32'd80: o_read_data = 32'd1303;
32'd84: o_read_data = 32'd38077715;
32'd88: o_read_data = 32'd1123875;
32'd92: o_read_data = 32'd4225757423;
32'd96: o_read_data = 32'd12656771;
32'd100: o_read_data = 32'd1303;
32'd104: o_read_data = 32'd33883411;
32'd108: o_read_data = 32'd16843027;
32'd112: o_read_data = 32'd4204785775;
32'd116: o_read_data = 32'd1819043144;
32'd120: o_read_data = 32'd1634934895;
32'd124: o_read_data = 32'd1919904873;
32'd128: o_read_data = 32'd2606;
32'd132: o_read_data = 32'd1952540759;
32'd136: o_read_data = 32'd1713402663;
32'd140: o_read_data = 32'd1646293615;
32'd144: o_read_data = 32'd1801545074;
32'd148: o_read_data = 32'd1953718630;
32'd152: o_read_data = 32'd2623;
default: o_read_data = 32'bX; // Default value
