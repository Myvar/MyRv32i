typedef enum reg [2:0] { 
PORT_ROM,
PORT_LRAM
} TargetPort;
