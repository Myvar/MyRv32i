`timescale 1ns / 1ps
`default_nettype none

module core #(
    parameter int AW = 32,
    parameter int DW = 32
) (
    input i_clk,
    input i_clk_en,
    input i_rst
);



endmodule
