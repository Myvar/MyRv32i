`ifndef OPCODE_SVH
`define OPCODE_SVH
typedef enum logic [8:0] {
  OP_NO_OP,
  OP_ADD,
  OP_SUB,
  OP_XOR,
  OP_OR,
  OP_AND,
  OP_SLL,
  OP_SRL,
  OP_SRA,
  OP_SLT,
  OP_SLTU,
  OP_ADDI,
  OP_XORI,
  OP_ORI,
  OP_ANDI,
  OP_SLLI,
  OP_SRLI,
  OP_SRAI,
  OP_SLTI,
  OP_SLTIU,
  OP_LB,
  OP_LH,
  OP_LW,
  OP_LBU,
  OP_LHU,
  OP_SB,
  OP_SH,
  OP_SW,
  OP_BEQ,
  OP_BNE,
  OP_BLT,
  OP_BGE,
  OP_BLTU,
  OP_BGEU,
  OP_JAL,
  OP_JALR,
  OP_LUI,
  OP_AUIPC,
  OP_ECALL,
  OP_EBREAK
} Opcode;

`endif  // MY_GUARD
