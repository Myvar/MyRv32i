32'd0: o_read_data = 32'd131;
default: o_read_data = 32'bX; // Default value
