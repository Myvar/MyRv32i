32'd0: o_read_data = 32'd131;
32'd4: o_read_data = 32'd605031459;
default: o_read_data = 32'bX; // Default value
